----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 12/18/2022 01:47:35 AM
-- Design Name: 
-- Module Name: dmux2_1 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity dmux2_1 is
Port (F:in std_logic_vector(63 downto 0);
      S:in std_logic;
      A,B:out std_logic_vector(63 downto 0));
end dmux2_1;

architecture Behavioral of dmux2_1 is
begin
process(F,S)
begin
  if S='0' then
    A<=F;
  else
    B<=F;
  end if;
end process;

end Behavioral;
